`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:55:47 06/24/2019 
// Design Name: 
// Module Name:    presetSR 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module presetSR(
    input pre,
    input clr,
    input clk,
    input s,
    input r,
    output q,
    output qb
    );


endmodule
