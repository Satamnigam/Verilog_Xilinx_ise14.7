`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   11:21:18 06/22/2019
// Design Name:   decod_3to8
// Module Name:   F:/my codes/decoder_3to8/decode_3_8.v
// Project Name:  decoder_3to8
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: decod_3to8
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module decode_3_8;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	decod_3to8 uut (
		.()
	);

	initial begin
		// Initialize Inputs
      i= 3'b010;
		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

